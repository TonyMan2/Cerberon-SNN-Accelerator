class pe_seq_item extends uvm_seq_item
    `uvm_component_utils(pe_seq_item)
    function new(string name = "pe_seq_item")
        
    endfunction